library verilog;
use verilog.vl_types.all;
entity testModule is
end testModule;
