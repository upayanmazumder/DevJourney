** Profile: "SCHEMATIC1-Max_power"  [ D:\upayanmazumder\DevJourney\Capture Cis Lite\Maximum Power Transfer Theorem\Maximum Power Transfer-PSpiceFiles\SCHEMATIC1\Max_power.sim ] 

** Creating circuit file "Max_power.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN PARAM RL 1 20 0.2 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
