** Profile: "SCHEMATIC1-RLC"  [ D:\upayanmazumder\DevJourney\Capture Cis Lite\Steady State Response of RLC Circuit\Steady State Response of RLC Circuit-PSpiceFiles\SCHEMATIC1\RLC.sim ] 

** Creating circuit file "RLC.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 100 0.1 100000
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
