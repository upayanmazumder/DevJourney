** Profile: "SCHEMATIC1-Half_Wave"  [ D:\upayanmazumder\DevJourney\Capture Cis Lite\Single Phase Rectifier\Half Wave Rectifier-PSpiceFiles\SCHEMATIC1\Half_Wave.sim ] 

** Creating circuit file "Half_Wave.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 0.04s 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
