library verilog;
use verilog.vl_types.all;
entity testModule2 is
end testModule2;
